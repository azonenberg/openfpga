localparam OP_TEST_RESET	=	3'h0;
localparam OP_RESET_IDLE	=	3'h1;
localparam OP_SELECT_IR		=	3'h2;
localparam OP_LEAVE_IR		=	3'h3;
localparam OP_SELECT_DR		=	3'h4;
localparam OP_LEAVE_DR		=	3'h5;
